`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.08.2019 03:22:17
// Design Name: 
// Module Name: to_ram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*

odule uart_rx_main(
    input logic uart_in_cable, reset, //reset con logica positiva
    input logic clock, //reloj de 100MHZ     IMPORTANTE!!!
    output logic [23:0] salida,
    output logic listo
*/

module to_ram(

    );
    
    uart
endmodule
